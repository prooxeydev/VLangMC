module io